// module Reset (output reg Reset, input GlobalReset);
//     always @( GlobalReset)
//     begin
//         if (GlobalReset == 1 )
//         Reset = 1;
//         else
//         Reset = 0;
//     end
// endmodule