//targetAddress Adder
module targetAddress(output [31:0] targetAddress_OUT, input[31:0] A, input[31:0] B);
     assign Adder_OUT = A + B;
endmodule
